`include "processor.v"

module processor_top;

endmodule