module shift();

endmodule